loader_inst : loader PORT MAP (
		noe_in	 => noe_in_sig
	);
